`timescale 1ns / 1ps

module ALUTestbench();
endmodule
